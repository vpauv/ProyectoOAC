library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory is
Port ( 
	dir : in STD_LOGIC_VECTOR (11 downto 0);
	data : out STD_LOGIC_VECTOR (97 downto 0));
end memory;

architecture Behavioral of memory is

begin
	process(dir)
	begin
	
		-- DATA FORMAT
		-- |    PRUEBA    |VF| Ins |                LIGA                 |
		--  P4 P3 P2 P1 P0 VF I1 I0 L11 L10 L9 L8 L7 L6 L5 L4 L3 L2 L1 L0 nCRI EB1 EB0 nWB EA1 EA0 nWA selbus UPA9 UPA8 UPA7 UPA6 UPA5 UPA4 UPA3 UPA2 UPA1 UPA0 nOEUPA nDUPA selmux nEX2 nEX1 nEX0 X2 X1 X0 EnaY nERA2 nERA1 nERA0 RA2 RA1 RA0 nEAP2 nEAP1 nEAP0 AP2 AP1 AP0 nEPC2 nEPC1 nEPC0 PC2 PC1 PC0 nCBD nAS nRW BD DINT HINT SET_IRQ SET_XIRQ B9 B8 B7 B6 B5 B4 B3 B2 B1 B0 CC CN CV CZ CI CH CX CS nHB ACCSEC

		-- Cadena por default: "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010"
		
		--if(dir=    X"000") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010";
		--elsif(dir= X"001") then data <= "00000" & "0" & "00" & "000000000000" & "00000000000000000000000000000000000000000000000000000000000000000000000000"; 
												  
		--FETCH			  
		if(dir=    X"000") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"001") then data <= "00000000000000000000000100100000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"002") then data <= "00000010000000000000100100100000000000110111000011100011100011100011111110000000000000000000000010";
		
		--LDAA(IMM)
		elsif(dir= X"860") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"861") then data <= "00000000000000000000100101000000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"862") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"863") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		--LDAB(IMM)
		elsif(dir= X"C60") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"C61") then data <= "00000000000000000000101000100000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"C62") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000100101000111000010";
		elsif(dir= X"C63") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		--ABA(INH)
		elsif(dir= X"1B0") then data <= "00000000000000000000111111100000000001111111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"1B1") then data <= "01111111000000000000100101000000000000000111000011100011100011100011111110000000000000001111010010";
		elsif(dir= X"1B2") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		--JMP(EXT)
		elsif(dir= X"7E0") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7E1") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir= X"7E2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7E3") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"7E4") then data <= "01111111000000000000100100100000000000110111000010000011100010010111111110000000000000000000000010";
		elsif(dir= X"7E5") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		--CPM(INH)
		elsif(dir= X"1C0") then data <= "00000000000000000000111111100000100001111111000011100011100011100011111110000000000000000000000011";
		elsif(dir= X"1C1") then data <= "01111111000000000000100100100000000000000111000011100011100011100011111110000000000000001111010010";
		elsif(dir= X"1C2") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
	
	   --JE(EXT)
		elsif(dir= X"7A0") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7A1") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir= X"7A2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"7A3") then data <= "00000001011110100101100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"7A4") then data <= "01111111000000000000100100100000000000110111000010000011100010010111111110000000000000000000000010";
		elsif(dir= X"7A5") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--JA(EXT)
		elsif(dir= X"6B0") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"6B1") then data <= "00000000000000000000100100100000000000110111000010110011100011100111111011000000000000000000000010";
		elsif(dir= X"6B2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"6B3") then data <= "10011101011010110101100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"6B4") then data <= "01111111000000000000100100100000000000110111000010000011100010010111111110000000000000000000000010";
		elsif(dir= X"6B5") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--LDX(IMM)
		elsif(dir= X"8D0") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"8D1") then data <= "00000000000000000000100100100000000000110110011011100011100011100111111010000000000000000000000010";
		elsif(dir= X"8D2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"8D3") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"8D4") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"8D5") then data <= "00000000000000000000100101000000000000110111000011100011100011100111111010000000000000000000000010";
		elsif(dir= X"8D6") then data <= "00000000000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"8D7") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--LDAA(DIR)
		elsif(dir= X"870") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"871") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir= X"872") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"873") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"874") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"875") then data <= "00000000000000000000100101000000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir= X"876") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"877") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--LDAB(DIR)
		elsif(dir= X"3C0") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir= X"3C1") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir= X"3C2") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir= X"3C3") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir= X"3C4") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir= X"3C5") then data <= "00000000000000000000101000100000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir= X"3C6") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir= X"3C7") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";

		--STAA(DIR)
		elsif(dir=X"A80") then data <= "00000000000000000000100111100001000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"A81") then data <= "00000000000000000000100100100000000000000111000010110011100011100011111110000000000000000000000010";
		elsif(dir=X"A82") then data <= "00000000000000000000100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir=X"A83") then data <= "00000000000000000000100100100000000000110111000011001111100011100111111010000000000000000000000010";
		elsif(dir=X"A84") then data <= "00000000000000000000100100100000000000110111000001100011100011100001111110000000000000000000000010";
		elsif(dir=X"A85") then data <= "00000000000000000000100101100000000000110111000011100011100011100011111000000000000000000000000010";
		elsif(dir=X"A86") then data <= "01111111000000000000100100100000000000110111000011100011100011100011111110000000010011000111000010";
		elsif(dir=X"A87") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		
		--MUL
		elsif(dir=X"F20") then data <= "00000000000000000000100111100000110000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F21") then data <= "00000000000000000000100100100011000010110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F22") then data <= "00000000000000000000100101000000001010000111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F23") then data <= "00001001111100101011100100100000000000100111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F24") then data <= "00000000000000000000111111100010000001110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F25") then data <= "00000000000000000000100100101010000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F26") then data <= "00000000000000000000100100101000000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F27") then data <= "01110001111100100011100101000000001011000111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F28") then data <= "00000000000000000000100100100010110010110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F29") then data <= "01111111000000000000101000100000000000000111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"F2A") then data <= "11000001000000000001100100100000000000110111000011100011100001100001111110000000000000000000000010";
		elsif(dir=X"F2B") then data <= "11000001111100100101100111100010000000110111000011100011100011100011111110000000000000000000000010";
		
		--EXTL
		elsif(dir=X"EA0") then data <= "00000000000000000000100100100101000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"EA1") then data <= "01111111000000000000101101000000000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"EA2") then data <= "11000001000000000001100100100000000000110111000011100011100011100011111110000000000000000000000010";
		
		
		--EXTH
		elsif(dir=X"EB0") then data <= "00000000000000000000100100100101000000110111000011100011100011100011111110000000000000000000000010";
		elsif(dir=X"EB1") then data <= "00000000000000000000100100100000000000110011000011100011100011100001111110000000000000000000000010";
		elsif(dir=X"EB2") then data <= "00000000000000000000110100100000000000110111000011100011100011100011111000000000000000000000000010";
		elsif(dir=X"EB3") then data <= "01111111000000000000100101000000000000110111000011100011100011100011111010000000000000000000000010";
		elsif(dir=X"EB4") then data <= "11000001000000000001100100100000000000110111000011100011100011100011111110000000000000000000000010";
		
		
		elsif(dir= X"200") then data <= "11000001000000000000100100100000000000110111000011100011100010010111011110000000000000000000000010";
		
		--else data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000000000000000000010"; -- Default
		----------------------------------------------
		
		
		
		----------------------------------------------
		
		else data <= "00000000000000000000100100100000000000110111000011100011100011100011111110000000000000000000000010";

		end if;
	end process;
end Behavioral;